module CLOCK_24(CLK, RESET, DEC, LED, SA, SW);
input CLK, RESET, DEC, SW;
output[7:0] LED;
output[3:0] SA;

wire[3:0] CNT10_SEC, CNT10_MIN, CNT10_HOUR, LED_TMP;
wire[2:0] CNT6_SEC, CNT6_MIN;
wire[1:0] CNT3_HOUR;
wire ENABLE, ENABLE_khz, MIN_CARRY,HOUR_CARRY,DAY_CARRY;
wire[7:0] LED_60;


ENABLE_GEN i0(.CLK(CLK), .RESET(RESET), .ENABLE(ENABLE), .ENABLE_khz(ENABLE_khz));
CNT60 i1(.CLK(CLK), .RESET(RESET), .DEC(DEC), .IN_CARRY(1'b1), .OUT_CARRY(MIN_CARRY), .ENABLE(ENABLE), .CNT10(CNT10_SEC), .CNT6(CNT6_SEC));
CNT60 i2(.CLK(CLK), .RESET(RESET), .DEC(DEC), .IN_CARRY(MIN_CARRY), .OUT_CARRY(HOUR_CARRY), .ENABLE(ENABLE), .CNT10(CNT10_MIN), .CNT6(CNT6_MIN));
CNT24 i3(.CLK(CLK), .RESET(RESET), .DEC(DEC), .IN_CARRY(HOUR_CARRY), .OUT_CARRY(DAY_CARRY), .ENABLE(ENABLE), .CNT10(CNT10_HOUR), .CNT3(CNT3_HOUR));
DCOUNT i4(.CLK(CLK), .ENABLE(ENABLE_khz), .L1(CNT10_SEC), .L2({1'b0,CNT6_SEC}), .L3(CNT10_MIN), .L4({1'b0,CNT6_MIN}), .L5(CNT10_HOUR), .L6({1'b0,1'b0,CNT3_HOUR}), .SA(SA), .L(LED_TMP), .SW(SW));
DECODER7 i5(.COUNT(LED_TMP), .LED(LED_60));

assign LED = ~LED_60;
endmodule